module tt_um_fpga_calculator (
    input  wire [7:0] ui_in,    // Dedicated inputs - connected to the input switches
    output wire [7:0] uo_out,   // Dedicated outputs - connected to the 7 segment display
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);


   wire reset = ! rst_n;

// ---------- Generated Code Inlined Here (before 1st \TLV) ----------
// Generated by SandPiper(TM) 1.14-2022/10/10-beta-Pro from Redwood EDA, LLC.
// (Installed here: /usr/local/mono/sandpiper/distro.)
// Redwood EDA, LLC does not claim intellectual property rights to this file and provides no warranty regarding its correctness or quality.


// For silencing unused signal messages.
`define BOGUS_USE(ignore)


genvar digit, input_label, leds, switch;


//
// Signals declared top-level.
//

// For $slideswitch.
logic [7:0] L0_slideswitch_a0;

// For $sseg_decimal_point_n.
logic L0_sseg_decimal_point_n_a0;

// For $sseg_digit_n.
logic [7:0] L0_sseg_digit_n_a0;

// For $sseg_segment_n.
logic [6:0] L0_sseg_segment_n_a0;

// For /fpga_pins/fpga|calc$diff.
logic [7:0] FpgaPins_Fpga_CALC_diff_a1,
            FpgaPins_Fpga_CALC_diff_a2;

// For /fpga_pins/fpga|calc$digit.
logic [3:0] FpgaPins_Fpga_CALC_digit_a3;

// For /fpga_pins/fpga|calc$mem.
logic [7:0] FpgaPins_Fpga_CALC_mem_a2,
            FpgaPins_Fpga_CALC_mem_a3,
            FpgaPins_Fpga_CALC_mem_a4;

// For /fpga_pins/fpga|calc$op.
logic [2:0] FpgaPins_Fpga_CALC_op_a0,
            FpgaPins_Fpga_CALC_op_a1,
            FpgaPins_Fpga_CALC_op_a2;

// For /fpga_pins/fpga|calc$out.
logic [7:0] FpgaPins_Fpga_CALC_out_a2,
            FpgaPins_Fpga_CALC_out_a3,
            FpgaPins_Fpga_CALC_out_a4;

// For /fpga_pins/fpga|calc$prod.
logic [7:0] FpgaPins_Fpga_CALC_prod_a1,
            FpgaPins_Fpga_CALC_prod_a2;

// For /fpga_pins/fpga|calc$quot.
logic [7:0] FpgaPins_Fpga_CALC_quot_a1,
            FpgaPins_Fpga_CALC_quot_a2;

// For /fpga_pins/fpga|calc$reset.
logic FpgaPins_Fpga_CALC_reset_a0,
      FpgaPins_Fpga_CALC_reset_a1,
      FpgaPins_Fpga_CALC_reset_a2;

// For /fpga_pins/fpga|calc$reset_or_valid.
logic FpgaPins_Fpga_CALC_reset_or_valid_a1,
      FpgaPins_Fpga_CALC_reset_or_valid_a2;

// For /fpga_pins/fpga|calc$sum.
logic [7:0] FpgaPins_Fpga_CALC_sum_a1,
            FpgaPins_Fpga_CALC_sum_a2;

// For /fpga_pins/fpga|calc$val1.
logic [7:0] FpgaPins_Fpga_CALC_val1_a1,
            FpgaPins_Fpga_CALC_val1_a2;

// For /fpga_pins/fpga|calc$val2.
logic [7:0] FpgaPins_Fpga_CALC_val2_a0,
            FpgaPins_Fpga_CALC_val2_a1;

// For /fpga_pins/fpga|calc$valid.
logic FpgaPins_Fpga_CALC_valid_a1,
      FpgaPins_Fpga_CALC_valid_a2;




   //
   // Scope: /fpga_pins
   //


      //
      // Scope: /fpga
      //


         //
         // Scope: |calc
         //

            // Staging of $diff.
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_diff_a2[7:0] <= FpgaPins_Fpga_CALC_diff_a1[7:0];

            // Staging of $mem.
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_mem_a3[7:0] <= FpgaPins_Fpga_CALC_mem_a2[7:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_mem_a4[7:0] <= FpgaPins_Fpga_CALC_mem_a3[7:0];

            // Staging of $op.
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_op_a1[2:0] <= FpgaPins_Fpga_CALC_op_a0[2:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_op_a2[2:0] <= FpgaPins_Fpga_CALC_op_a1[2:0];

            // Staging of $out.
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_out_a3[7:0] <= FpgaPins_Fpga_CALC_out_a2[7:0];
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_out_a4[7:0] <= FpgaPins_Fpga_CALC_out_a3[7:0];

            // Staging of $prod.
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_prod_a2[7:0] <= FpgaPins_Fpga_CALC_prod_a1[7:0];

            // Staging of $quot.
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_quot_a2[7:0] <= FpgaPins_Fpga_CALC_quot_a1[7:0];

            // Staging of $reset.
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_reset_a1 <= FpgaPins_Fpga_CALC_reset_a0;
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_reset_a2 <= FpgaPins_Fpga_CALC_reset_a1;

            // Staging of $reset_or_valid.
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_reset_or_valid_a2 <= FpgaPins_Fpga_CALC_reset_or_valid_a1;

            // Staging of $sum.
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_sum_a2[7:0] <= FpgaPins_Fpga_CALC_sum_a1[7:0];

            // Staging of $val1.
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_val1_a2[7:0] <= FpgaPins_Fpga_CALC_val1_a1[7:0];

            // Staging of $val2.
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_val2_a1[7:0] <= FpgaPins_Fpga_CALC_val2_a0[7:0];

            // Staging of $valid.
            always_ff @(posedge clk) FpgaPins_Fpga_CALC_valid_a2 <= FpgaPins_Fpga_CALC_valid_a1;




// ---------- Generated Code Ends ----------
//_\TLV
   /* verilator lint_off UNOPTFLAT */
   // Connect Tiny Tapeout I/Os to Virtual FPGA Lab.
   //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/af18805ea79802b83477cf86aff503e97ed7394a/tlvlib/tinytapeoutlib.tlv 67   // Instantiated from top.tlv, 859 as: m5+tt_connections()
      assign L0_slideswitch_a0[7:0] = ui_in;
      assign L0_sseg_segment_n_a0[6:0] = uo_out[6:0];
      assign L0_sseg_decimal_point_n_a0 = uo_out[7];
      assign L0_sseg_digit_n_a0[7:0] = 8'b11111110;
   //_\end_source

   // Instantiate the Virtual FPGA Lab.
   //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv 307   // Instantiated from top.tlv, 862 as: m5+board(/top, /fpga, 7, $, , hidden_solution)

      //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv 355   // Instantiated from /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv, 309 as: m4+thanks(m5__l(309)m5_eval(m5_get(BOARD_THANKS_ARGS)))
         //_/thanks

      //_\end_source


      // Board VIZ.

      // Board Image.

      //_/fpga_pins

         //_/fpga
            //_\source top.tlv 205   // Instantiated from /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv, 340 as: m4+hidden_solution.
               //_\source top.tlv 208   // Instantiated from top.tlv, 206 as: m5+call(m5__l(206)m5_call(if,m5_get(CalcLab), calc_solution, cpu_solution))
                  /* verilator lint_off WIDTH */
                  //_|calc

                     // ============================================================================================================


                     //_@0
                        assign FpgaPins_Fpga_CALC_reset_a0 = reset;

                     //_@0
                        // Board inputs
                        assign FpgaPins_Fpga_CALC_op_a0[2:0] = ui_in[7:5];
                        assign FpgaPins_Fpga_CALC_val2_a0[7:0] = {3'b0, ui_in[4:0]};

                     //_@1

                        //$reset = *reset;
                        assign FpgaPins_Fpga_CALC_val1_a1[7:0] = FpgaPins_Fpga_CALC_out_a3;


                        assign FpgaPins_Fpga_CALC_valid_a1 = FpgaPins_Fpga_CALC_reset_a1 ? 1'b0 : FpgaPins_Fpga_CALC_valid_a2 + 1'b1;
                        assign FpgaPins_Fpga_CALC_reset_or_valid_a1 = FpgaPins_Fpga_CALC_valid_a1 || FpgaPins_Fpga_CALC_reset_a1;













                     //_?$reset_or_valid
                        //_@1
                           assign FpgaPins_Fpga_CALC_sum_a1[7:0] = FpgaPins_Fpga_CALC_val1_a1 + FpgaPins_Fpga_CALC_val2_a1;
                           assign FpgaPins_Fpga_CALC_diff_a1[7:0] = FpgaPins_Fpga_CALC_val1_a1 - FpgaPins_Fpga_CALC_val2_a1;
                           assign FpgaPins_Fpga_CALC_prod_a1[7:0] = FpgaPins_Fpga_CALC_val1_a1 + FpgaPins_Fpga_CALC_val2_a1;
                           assign FpgaPins_Fpga_CALC_quot_a1[7:0] = FpgaPins_Fpga_CALC_val1_a1 - FpgaPins_Fpga_CALC_val2_a1;
                        //_@2

                           assign FpgaPins_Fpga_CALC_mem_a2[7:0] = FpgaPins_Fpga_CALC_reset_a2           ? 8'b0 :
                                           (FpgaPins_Fpga_CALC_op_a2[2:0] == 3'b101) ? FpgaPins_Fpga_CALC_val1_a2 :
                                                              FpgaPins_Fpga_CALC_mem_a4;

                           assign FpgaPins_Fpga_CALC_out_a2[7:0] = FpgaPins_Fpga_CALC_reset_a2           ? 8'b0 :
                                        (FpgaPins_Fpga_CALC_op_a2 == 3'b000) ? FpgaPins_Fpga_CALC_sum_a2  :
                                        (FpgaPins_Fpga_CALC_op_a2 == 3'b001) ? FpgaPins_Fpga_CALC_diff_a2 :
                                        (FpgaPins_Fpga_CALC_op_a2 == 3'b010) ? FpgaPins_Fpga_CALC_prod_a2 :
                                        (FpgaPins_Fpga_CALC_op_a2 == 3'b011) ? FpgaPins_Fpga_CALC_quot_a2 :
                                        (FpgaPins_Fpga_CALC_op_a2 == 3'b100) ? FpgaPins_Fpga_CALC_mem_a4 : FpgaPins_Fpga_CALC_out_a4;


















                     //_@3
                        assign FpgaPins_Fpga_CALC_digit_a3[3:0] = FpgaPins_Fpga_CALC_out_a3[3:0];
                        assign uo_out =
                           FpgaPins_Fpga_CALC_digit_a3 == 4'h0 ? 8'b11000000 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'h1 ? 8'b11111001 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'h2 ? 8'b10100100 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'h3 ? 8'b10110000 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'h4 ? 8'b10011001 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'h5 ? 8'b10010010 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'h6 ? 8'b10000010 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'h7 ? 8'b11111000 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'h8 ? 8'b10000000 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'h9 ? 8'b10010000 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'hA ? 8'b10001000 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'hB ? 8'b10000011 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'hC ? 8'b11000110 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'hD ? 8'b10100001 :
                           FpgaPins_Fpga_CALC_digit_a3 == 4'hE ? 8'b10000110 :
                                            8'b10001110;





                  // ============================================================================================================

                  // Connect Tiny Tapeout outputs.
                  // (*uo_out connected above.)
                  // assign uio_out = 8'b0;
                  // assign uio_oe = 8'b0;
               //_\end_source

            //_\end_source

      // LEDs.


      // 7-Segment
      //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv 395   // Instantiated from /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv, 346 as: m4+fpga_sseg.
         for (digit = 0; digit <= 0; digit++) begin : L1_Digit //_/digit

            for (leds = 0; leds <= 7; leds++) begin : L2_Leds //_/leds

               // For $viz_lit.
               logic L2_viz_lit_a0;

               assign L2_viz_lit_a0 = (! L0_sseg_digit_n_a0[digit]) && ! ((leds == 7) ? L0_sseg_decimal_point_n_a0 : L0_sseg_segment_n_a0[leds % 7]);

            end
         end
      //_\end_source

      // slideswitches
      //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv 454   // Instantiated from /raw.githubusercontent.com/osfpga/VirtualFPGALab/a069f1e4e19adc829b53237b3e0b5d6763dc3194/tlvlib/fpgaincludes.tlv, 349 as: m4+fpga_switch.
         for (switch = 0; switch <= 7; switch++) begin : L1_Switch //_/switch

            // For $viz_switch.
            logic L1_viz_switch_a0;

            assign L1_viz_switch_a0 = L0_slideswitch_a0[switch];

         end
      //_\end_source

      // pushbuttons

   //_\end_source
   // Label the switch inputs [0..7] (1..8 on the physical switch panel) (bottom-to-top).
   //_\source /raw.githubusercontent.com/osfpga/VirtualFPGALab/af18805ea79802b83477cf86aff503e97ed7394a/tlvlib/tinytapeoutlib.tlv 73   // Instantiated from top.tlv, 864 as: m5+tt_input_labels_viz(m5_get(input_labels))
      for (input_label = 0; input_label <= 7; input_label++) begin : L1_InputLabel //_/input_label

      end
   //_\end_source

//_\SV
endmodule


// Undefine macros defined by SandPiper.
`undef BOGUS_USE
